module vk

import misc

pub struct Mesh {
pub:
	verticies []misc.Vertex
	indicies  []u32
}
