module vulkan

#flag -L @VMODROOT/libs/vulkan/libvulkan.so
#flag -lvulkan
#flag -I @VMODROOT/libs/vulkan/latest/x86_64/include
#include "vulkan/vulkan.h"
