module vulkan

fn C.VK_MAKE_VERSION(u32, u32, u32) u32
