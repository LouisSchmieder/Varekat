module glfw

#pkgconfig glfw3
#include <GLFW/glfw3.h>
