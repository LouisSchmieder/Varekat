module vulkan

pub enum ShaderType {
	fragment = 0x00000010
	vertex = 0x00000001
}

pub enum AttachmentLoadOp {
	vk_attachment_load_op_load = 0
	vk_attachment_load_op_clear = 1
	vk_attachment_load_op_dont_care = 2
}

pub enum AttachmentStoreOp {
	vk_attachment_store_op_store = 0
	vk_attachment_store_op_dont_care = 1
	vk_attachment_store_op_none_ext = 1000301000
}

pub enum ImageLayout {
	vk_image_layout_undefined = 0
	vk_image_layout_general = 1
	vk_image_layout_color_attachment_optimal = 2
	vk_image_layout_depth_stencil_attachment_optimal = 3
	vk_image_layout_depth_stencil_read_only_optimal = 4
	vk_image_layout_shader_read_only_optimal = 5
	vk_image_layout_transfer_src_optimal = 6
	vk_image_layout_transfer_dst_optimal = 7
	vk_image_layout_preinitialized = 8
	vk_image_layout_depth_read_only_stencil_attachment_optimal = 1000117000
	vk_image_layout_depth_attachment_stencil_read_only_optimal = 1000117001
	vk_image_layout_depth_attachment_optimal = 1000241000
	vk_image_layout_depth_read_only_optimal = 1000241001
	vk_image_layout_stencil_attachment_optimal = 1000241002
	vk_image_layout_stencil_read_only_optimal = 1000241003
	vk_image_layout_present_src_khr = 1000001002
	vk_image_layout_video_decode_dst_khr = 1000024000
	vk_image_layout_video_decode_src_khr = 1000024001
	vk_image_layout_video_decode_dpb_khr = 1000024002
	vk_image_layout_shared_present_khr = 1000111000
	vk_image_layout_fragment_density_map_optimal_ext = 1000218000
	vk_image_layout_fragment_shading_rate_attachment_optimal_khr = 1000164003
	vk_image_layout_video_encode_dst_khr = 1000299000
	vk_image_layout_video_encode_src_khr = 1000299001
	vk_image_layout_video_encode_dpb_khr = 1000299002
	vk_image_layout_read_only_optimal_khr = 1000314000
	vk_image_layout_attachment_optimal_khr = 1000314001
}

pub enum LogicOp {
	vk_logic_op_clear = 0
	vk_logic_op_and = 1
	vk_logic_op_and_reverse = 2
	vk_logic_op_copy = 3
	vk_logic_op_and_inverted = 4
	vk_logic_op_no_op = 5
	vk_logic_op_xor = 6
	vk_logic_op_or = 7
	vk_logic_op_nor = 8
	vk_logic_op_equivalent = 9
	vk_logic_op_invert = 10
	vk_logic_op_or_reverse = 11
	vk_logic_op_copy_inverted = 12
	vk_logic_op_or_inverted = 13
	vk_logic_op_nand = 14
	vk_logic_op_set = 15
	vk_logic_op_max_enum = 0x7fffffff
}

pub enum BlendFactor {
	vk_blend_factor_zero = 0
	vk_blend_factor_one = 1
	vk_blend_factor_src_color = 2
	vk_blend_factor_one_minus_src_color = 3
	vk_blend_factor_dst_color = 4
	vk_blend_factor_one_minus_dst_color = 5
	vk_blend_factor_src_alpha = 6
	vk_blend_factor_one_minus_src_alpha = 7
	vk_blend_factor_dst_alpha = 8
	vk_blend_factor_one_minus_dst_alpha = 9
	vk_blend_factor_constant_color = 10
	vk_blend_factor_one_minus_constant_color = 11
	vk_blend_factor_constant_alpha = 12
	vk_blend_factor_one_minus_constant_alpha = 13
	vk_blend_factor_src_alpha_saturate = 14
	vk_blend_factor_src1_color = 15
	vk_blend_factor_one_minus_src1_color = 16
	vk_blend_factor_src1_alpha = 17
	vk_blend_factor_one_minus_src1_alpha = 18
	vk_blend_factor_max_enum = 0x7fffffff
}

pub enum BlendOp {
	vk_blend_op_add = 0
	vk_blend_op_subtract = 1
	vk_blend_op_reverse_subtract = 2
	vk_blend_op_min = 3
	vk_blend_op_max = 4
	vk_blend_op_zero_ext = 1000148000
	vk_blend_op_src_ext = 1000148001
	vk_blend_op_dst_ext = 1000148002
	vk_blend_op_src_over_ext = 1000148003
	vk_blend_op_dst_over_ext = 1000148004
	vk_blend_op_src_in_ext = 1000148005
	vk_blend_op_dst_in_ext = 1000148006
	vk_blend_op_src_out_ext = 1000148007
	vk_blend_op_dst_out_ext = 1000148008
	vk_blend_op_src_atop_ext = 1000148009
	vk_blend_op_dst_atop_ext = 1000148010
	vk_blend_op_xor_ext = 1000148011
	vk_blend_op_multiply_ext = 1000148012
	vk_blend_op_screen_ext = 1000148013
	vk_blend_op_overlay_ext = 1000148014
	vk_blend_op_darken_ext = 1000148015
	vk_blend_op_lighten_ext = 1000148016
	vk_blend_op_colordodge_ext = 1000148017
	vk_blend_op_colorburn_ext = 1000148018
	vk_blend_op_hardlight_ext = 1000148019
	vk_blend_op_softlight_ext = 1000148020
	vk_blend_op_difference_ext = 1000148021
	vk_blend_op_exclusion_ext = 1000148022
	vk_blend_op_invert_ext = 1000148023
	vk_blend_op_invert_rgb_ext = 1000148024
	vk_blend_op_lineardodge_ext = 1000148025
	vk_blend_op_linearburn_ext = 1000148026
	vk_blend_op_vividlight_ext = 1000148027
	vk_blend_op_linearlight_ext = 1000148028
	vk_blend_op_pinlight_ext = 1000148029
	vk_blend_op_hardmix_ext = 1000148030
	vk_blend_op_hsl_hue_ext = 1000148031
	vk_blend_op_hsl_saturation_ext = 1000148032
	vk_blend_op_hsl_color_ext = 1000148033
	vk_blend_op_hsl_luminosity_ext = 1000148034
	vk_blend_op_plus_ext = 1000148035
	vk_blend_op_plus_clamped_ext = 1000148036
	vk_blend_op_plus_clamped_alpha_ext = 1000148037
	vk_blend_op_plus_darker_ext = 1000148038
	vk_blend_op_minus_ext = 1000148039
	vk_blend_op_minus_clamped_ext = 1000148040
	vk_blend_op_contrast_ext = 1000148041
	vk_blend_op_invert_ovg_ext = 1000148042
	vk_blend_op_red_ext = 1000148043
	vk_blend_op_green_ext = 1000148044
	vk_blend_op_blue_ext = 1000148045
	vk_blend_op_max_enum = 0x7fffffff
}

pub enum StructureType {
	vk_structure_type_application_info = 0
	vk_structure_type_instance_create_info = 1
	vk_structure_type_device_queue_create_info = 2
	vk_structure_type_device_create_info = 3
	vk_structure_type_submit_info = 4
	vk_structure_type_memory_allocate_info = 5
	vk_structure_type_mapped_memory_range = 6
	vk_structure_type_bind_sparse_info = 7
	vk_structure_type_fence_create_info = 8
	vk_structure_type_semaphore_create_info = 9
	vk_structure_type_event_create_info = 10
	vk_structure_type_query_pool_create_info = 11
	vk_structure_type_buffer_create_info = 12
	vk_structure_type_buffer_view_create_info = 13
	vk_structure_type_image_create_info = 14
	vk_structure_type_image_view_create_info = 15
	vk_structure_type_shader_module_create_info = 16
	vk_structure_type_pipeline_cache_create_info = 17
	vk_structure_type_pipeline_shader_stage_create_info = 18
	vk_structure_type_pipeline_vertex_input_state_create_info = 19
	vk_structure_type_pipeline_input_assembly_state_create_info = 20
	vk_structure_type_pipeline_tessellation_state_create_info = 21
	vk_structure_type_pipeline_viewport_state_create_info = 22
	vk_structure_type_pipeline_rasterization_state_create_info = 23
	vk_structure_type_pipeline_multisample_state_create_info = 24
	vk_structure_type_pipeline_depth_stencil_state_create_info = 25
	vk_structure_type_pipeline_color_blend_state_create_info = 26
	vk_structure_type_pipeline_dynamic_state_create_info = 27
	vk_structure_type_graphics_pipeline_create_info = 28
	vk_structure_type_compute_pipeline_create_info = 29
	vk_structure_type_pipeline_layout_create_info = 30
	vk_structure_type_sampler_create_info = 31
	vk_structure_type_descriptor_set_layout_create_info = 32
	vk_structure_type_descriptor_pool_create_info = 33
	vk_structure_type_descriptor_set_allocate_info = 34
	vk_structure_type_write_descriptor_set = 35
	vk_structure_type_copy_descriptor_set = 36
	vk_structure_type_framebuffer_create_info = 37
	vk_structure_type_render_pass_create_info = 38
	vk_structure_type_command_pool_create_info = 39
	vk_structure_type_command_buffer_allocate_info = 40
	vk_structure_type_command_buffer_inheritance_info = 41
	vk_structure_type_command_buffer_begin_info = 42
	vk_structure_type_render_pass_begin_info = 43
	vk_structure_type_buffer_memory_barrier = 44
	vk_structure_type_image_memory_barrier = 45
	vk_structure_type_memory_barrier = 46
	vk_structure_type_loader_instance_create_info = 47
	vk_structure_type_loader_device_create_info = 48
	vk_structure_type_physical_device_subgroup_properties = 1000094000
	vk_structure_type_bind_buffer_memory_info = 1000157000
	vk_structure_type_bind_image_memory_info = 1000157001
	vk_structure_type_physical_device_16bit_storage_features = 1000083000
	vk_structure_type_memory_dedicated_requirements = 1000127000
	vk_structure_type_memory_dedicated_allocate_info = 1000127001
	vk_structure_type_memory_allocate_flags_info = 1000060000
	vk_structure_type_device_group_render_pass_begin_info = 1000060003
	vk_structure_type_device_group_command_buffer_begin_info = 1000060004
	vk_structure_type_device_group_submit_info = 1000060005
	vk_structure_type_device_group_bind_sparse_info = 1000060006
	vk_structure_type_bind_buffer_memory_device_group_info = 1000060013
	vk_structure_type_bind_image_memory_device_group_info = 1000060014
	vk_structure_type_physical_device_group_properties = 1000070000
	vk_structure_type_device_group_device_create_info = 1000070001
	vk_structure_type_buffer_memory_requirements_info_2 = 1000146000
	vk_structure_type_image_memory_requirements_info_2 = 1000146001
	vk_structure_type_image_sparse_memory_requirements_info_2 = 1000146002
	vk_structure_type_memory_requirements_2 = 1000146003
	vk_structure_type_sparse_image_memory_requirements_2 = 1000146004
	vk_structure_type_physical_device_features_2 = 1000059000
	vk_structure_type_physical_device_properties_2 = 1000059001
	vk_structure_type_format_properties_2 = 1000059002
	vk_structure_type_image_format_properties_2 = 1000059003
	vk_structure_type_physical_device_image_format_info_2 = 1000059004
	vk_structure_type_queue_family_properties_2 = 1000059005
	vk_structure_type_physical_device_memory_properties_2 = 1000059006
	vk_structure_type_sparse_image_format_properties_2 = 1000059007
	vk_structure_type_physical_device_sparse_image_format_info_2 = 1000059008
	vk_structure_type_physical_device_point_clipping_properties = 1000117000
	vk_structure_type_render_pass_input_attachment_aspect_create_info = 1000117001
	vk_structure_type_image_view_usage_create_info = 1000117002
	vk_structure_type_pipeline_tessellation_domain_origin_state_create_info = 1000117003
	vk_structure_type_render_pass_multiview_create_info = 1000053000
	vk_structure_type_physical_device_multiview_features = 1000053001
	vk_structure_type_physical_device_multiview_properties = 1000053002
	vk_structure_type_physical_device_variable_pointers_features = 1000120000
	vk_structure_type_protected_submit_info = 1000145000
	vk_structure_type_physical_device_protected_memory_features = 1000145001
	vk_structure_type_physical_device_protected_memory_properties = 1000145002
	vk_structure_type_device_queue_info_2 = 1000145003
	vk_structure_type_sampler_ycbcr_conversion_create_info = 1000156000
	vk_structure_type_sampler_ycbcr_conversion_info = 1000156001
	vk_structure_type_bind_image_plane_memory_info = 1000156002
	vk_structure_type_image_plane_memory_requirements_info = 1000156003
	vk_structure_type_physical_device_sampler_ycbcr_conversion_features = 1000156004
	vk_structure_type_sampler_ycbcr_conversion_image_format_properties = 1000156005
	vk_structure_type_descriptor_update_template_create_info = 1000085000
	vk_structure_type_physical_device_external_image_format_info = 1000071000
	vk_structure_type_external_image_format_properties = 1000071001
	vk_structure_type_physical_device_external_buffer_info = 1000071002
	vk_structure_type_external_buffer_properties = 1000071003
	vk_structure_type_physical_device_id_properties = 1000071004
	vk_structure_type_external_memory_buffer_create_info = 1000072000
	vk_structure_type_external_memory_image_create_info = 1000072001
	vk_structure_type_export_memory_allocate_info = 1000072002
	vk_structure_type_physical_device_external_fence_info = 1000112000
	vk_structure_type_external_fence_properties = 1000112001
	vk_structure_type_export_fence_create_info = 1000113000
	vk_structure_type_export_semaphore_create_info = 1000077000
	vk_structure_type_physical_device_external_semaphore_info = 1000076000
	vk_structure_type_external_semaphore_properties = 1000076001
	vk_structure_type_physical_device_maintenance_3_properties = 1000168000
	vk_structure_type_descriptor_set_layout_support = 1000168001
	vk_structure_type_physical_device_shader_draw_parameters_features = 1000063000
	vk_structure_type_physical_device_vulkan_1_1_features = 49
	vk_structure_type_physical_device_vulkan_1_1_properties = 50
	vk_structure_type_physical_device_vulkan_1_2_features = 51
	vk_structure_type_physical_device_vulkan_1_2_properties = 52
	vk_structure_type_image_format_list_create_info = 1000147000
	vk_structure_type_attachment_description_2 = 1000109000
	vk_structure_type_attachment_reference_2 = 1000109001
	vk_structure_type_subpass_description_2 = 1000109002
	vk_structure_type_subpass_dependency_2 = 1000109003
	vk_structure_type_render_pass_create_info_2 = 1000109004
	vk_structure_type_subpass_begin_info = 1000109005
	vk_structure_type_subpass_end_info = 1000109006
	vk_structure_type_physical_device_8bit_storage_features = 1000177000
	vk_structure_type_physical_device_driver_properties = 1000196000
	vk_structure_type_physical_device_shader_atomic_int64_features = 1000180000
	vk_structure_type_physical_device_shader_float16_int8_features = 1000082000
	vk_structure_type_physical_device_float_controls_properties = 1000197000
	vk_structure_type_descriptor_set_layout_binding_flags_create_info = 1000161000
	vk_structure_type_physical_device_descriptor_indexing_features = 1000161001
	vk_structure_type_physical_device_descriptor_indexing_properties = 1000161002
	vk_structure_type_descriptor_set_variable_descriptor_count_allocate_info = 1000161003
	vk_structure_type_descriptor_set_variable_descriptor_count_layout_support = 1000161004
	vk_structure_type_physical_device_depth_stencil_resolve_properties = 1000199000
	vk_structure_type_subpass_description_depth_stencil_resolve = 1000199001
	vk_structure_type_physical_device_scalar_block_layout_features = 1000221000
	vk_structure_type_image_stencil_usage_create_info = 1000246000
	vk_structure_type_physical_device_sampler_filter_minmax_properties = 1000130000
	vk_structure_type_sampler_reduction_mode_create_info = 1000130001
	vk_structure_type_physical_device_vulkan_memory_model_features = 1000211000
	vk_structure_type_physical_device_imageless_framebuffer_features = 1000108000
	vk_structure_type_framebuffer_attachments_create_info = 1000108001
	vk_structure_type_framebuffer_attachment_image_info = 1000108002
	vk_structure_type_render_pass_attachment_begin_info = 1000108003
	vk_structure_type_physical_device_uniform_buffer_standard_layout_features = 1000253000
	vk_structure_type_physical_device_shader_subgroup_extended_types_features = 1000175000
	vk_structure_type_physical_device_separate_depth_stencil_layouts_features = 1000241000
	vk_structure_type_attachment_reference_stencil_layout = 1000241001
	vk_structure_type_attachment_description_stencil_layout = 1000241002
	vk_structure_type_physical_device_host_query_reset_features = 1000261000
	vk_structure_type_physical_device_timeline_semaphore_features = 1000207000
	vk_structure_type_physical_device_timeline_semaphore_properties = 1000207001
	vk_structure_type_semaphore_type_create_info = 1000207002
	vk_structure_type_timeline_semaphore_submit_info = 1000207003
	vk_structure_type_semaphore_wait_info = 1000207004
	vk_structure_type_semaphore_signal_info = 1000207005
	vk_structure_type_physical_device_buffer_device_address_features = 1000257000
	vk_structure_type_buffer_device_address_info = 1000244001
	vk_structure_type_buffer_opaque_capture_address_create_info = 1000257002
	vk_structure_type_memory_opaque_capture_address_allocate_info = 1000257003
	vk_structure_type_device_memory_opaque_capture_address_info = 1000257004
	vk_structure_type_swapchain_create_info_khr = 1000001000
	vk_structure_type_present_info_khr = 1000001001
	vk_structure_type_device_group_present_capabilities_khr = 1000060007
	vk_structure_type_image_swapchain_create_info_khr = 1000060008
	vk_structure_type_bind_image_memory_swapchain_info_khr = 1000060009
	vk_structure_type_acquire_next_image_info_khr = 1000060010
	vk_structure_type_device_group_present_info_khr = 1000060011
	vk_structure_type_device_group_swapchain_create_info_khr = 1000060012
	vk_structure_type_display_mode_create_info_khr = 1000002000
	vk_structure_type_display_surface_create_info_khr = 1000002001
	vk_structure_type_display_present_info_khr = 1000003000
	vk_structure_type_xlib_surface_create_info_khr = 1000004000
	vk_structure_type_xcb_surface_create_info_khr = 1000005000
	vk_structure_type_wayland_surface_create_info_khr = 1000006000
	vk_structure_type_android_surface_create_info_khr = 1000008000
	vk_structure_type_win32_surface_create_info_khr = 1000009000
	vk_structure_type_debug_report_callback_create_info_ext = 1000011000
	vk_structure_type_pipeline_rasterization_state_rasterization_order_amd = 1000018000
	vk_structure_type_debug_marker_object_name_info_ext = 1000022000
	vk_structure_type_debug_marker_object_tag_info_ext = 1000022001
	vk_structure_type_debug_marker_marker_info_ext = 1000022002
	vk_structure_type_video_profile_khr = 1000023000
	vk_structure_type_video_capabilities_khr = 1000023001
	vk_structure_type_video_picture_resource_khr = 1000023002
	vk_structure_type_video_get_memory_properties_khr = 1000023003
	vk_structure_type_video_bind_memory_khr = 1000023004
	vk_structure_type_video_session_create_info_khr = 1000023005
	vk_structure_type_video_session_parameters_create_info_khr = 1000023006
	vk_structure_type_video_session_parameters_update_info_khr = 1000023007
	vk_structure_type_video_begin_coding_info_khr = 1000023008
	vk_structure_type_video_end_coding_info_khr = 1000023009
	vk_structure_type_video_coding_control_info_khr = 1000023010
	vk_structure_type_video_reference_slot_khr = 1000023011
	vk_structure_type_video_queue_family_properties_2_khr = 1000023012
	vk_structure_type_video_profiles_khr = 1000023013
	vk_structure_type_physical_device_video_format_info_khr = 1000023014
	vk_structure_type_video_format_properties_khr = 1000023015
	vk_structure_type_video_decode_info_khr = 1000024000
	vk_structure_type_dedicated_allocation_image_create_info_nv = 1000026000
	vk_structure_type_dedicated_allocation_buffer_create_info_nv = 1000026001
	vk_structure_type_dedicated_allocation_memory_allocate_info_nv = 1000026002
	vk_structure_type_physical_device_transform_feedback_features_ext = 1000028000
	vk_structure_type_physical_device_transform_feedback_properties_ext = 1000028001
	vk_structure_type_pipeline_rasterization_state_stream_create_info_ext = 1000028002
	vk_structure_type_cu_module_create_info_nvx = 1000029000
	vk_structure_type_cu_function_create_info_nvx = 1000029001
	vk_structure_type_cu_launch_info_nvx = 1000029002
	vk_structure_type_image_view_handle_info_nvx = 1000030000
	vk_structure_type_image_view_address_properties_nvx = 1000030001
	vk_structure_type_video_encode_h264_capabilities_ext = 1000038000
	vk_structure_type_video_encode_h264_session_create_info_ext = 1000038001
	vk_structure_type_video_encode_h264_session_parameters_create_info_ext = 1000038002
	vk_structure_type_video_encode_h264_session_parameters_add_info_ext = 1000038003
	vk_structure_type_video_encode_h264_vcl_frame_info_ext = 1000038004
	vk_structure_type_video_encode_h264_dpb_slot_info_ext = 1000038005
	vk_structure_type_video_encode_h264_nalu_slice_ext = 1000038006
	vk_structure_type_video_encode_h264_emit_picture_parameters_ext = 1000038007
	vk_structure_type_video_encode_h264_profile_ext = 1000038008
	vk_structure_type_video_decode_h264_capabilities_ext = 1000040000
	vk_structure_type_video_decode_h264_session_create_info_ext = 1000040001
	vk_structure_type_video_decode_h264_picture_info_ext = 1000040002
	vk_structure_type_video_decode_h264_mvc_ext = 1000040003
	vk_structure_type_video_decode_h264_profile_ext = 1000040004
	vk_structure_type_video_decode_h264_session_parameters_create_info_ext = 1000040005
	vk_structure_type_video_decode_h264_session_parameters_add_info_ext = 1000040006
	vk_structure_type_video_decode_h264_dpb_slot_info_ext = 1000040007
	vk_structure_type_texture_lod_gather_format_properties_amd = 1000041000
	vk_structure_type_stream_descriptor_surface_create_info_ggp = 1000049000
	vk_structure_type_physical_device_corner_sampled_image_features_nv = 1000050000
	vk_structure_type_external_memory_image_create_info_nv = 1000056000
	vk_structure_type_export_memory_allocate_info_nv = 1000056001
	vk_structure_type_import_memory_win32_handle_info_nv = 1000057000
	vk_structure_type_export_memory_win32_handle_info_nv = 1000057001
	vk_structure_type_win32_keyed_mutex_acquire_release_info_nv = 1000058000
	vk_structure_type_validation_flags_ext = 1000061000
	vk_structure_type_vi_surface_create_info_nn = 1000062000
	vk_structure_type_physical_device_texture_compression_astc_hdr_features_ext = 1000066000
	vk_structure_type_image_view_astc_decode_mode_ext = 1000067000
	vk_structure_type_physical_device_astc_decode_features_ext = 1000067001
	vk_structure_type_import_memory_win32_handle_info_khr = 1000073000
	vk_structure_type_export_memory_win32_handle_info_khr = 1000073001
	vk_structure_type_memory_win32_handle_properties_khr = 1000073002
	vk_structure_type_memory_get_win32_handle_info_khr = 1000073003
	vk_structure_type_import_memory_fd_info_khr = 1000074000
	vk_structure_type_memory_fd_properties_khr = 1000074001
	vk_structure_type_memory_get_fd_info_khr = 1000074002
	vk_structure_type_win32_keyed_mutex_acquire_release_info_khr = 1000075000
	vk_structure_type_import_semaphore_win32_handle_info_khr = 1000078000
	vk_structure_type_export_semaphore_win32_handle_info_khr = 1000078001
	vk_structure_type_d3d12_fence_submit_info_khr = 1000078002
	vk_structure_type_semaphore_get_win32_handle_info_khr = 1000078003
	vk_structure_type_import_semaphore_fd_info_khr = 1000079000
	vk_structure_type_semaphore_get_fd_info_khr = 1000079001
	vk_structure_type_physical_device_push_descriptor_properties_khr = 1000080000
	vk_structure_type_command_buffer_inheritance_conditional_rendering_info_ext = 1000081000
	vk_structure_type_physical_device_conditional_rendering_features_ext = 1000081001
	vk_structure_type_conditional_rendering_begin_info_ext = 1000081002
	vk_structure_type_present_regions_khr = 1000084000
	vk_structure_type_pipeline_viewport_w_scaling_state_create_info_nv = 1000087000
	vk_structure_type_surface_capabilities_2_ext = 1000090000
	vk_structure_type_display_power_info_ext = 1000091000
	vk_structure_type_device_event_info_ext = 1000091001
	vk_structure_type_display_event_info_ext = 1000091002
	vk_structure_type_swapchain_counter_create_info_ext = 1000091003
	vk_structure_type_present_times_info_google = 1000092000
	vk_structure_type_physical_device_multiview_per_view_attributes_properties_nvx = 1000097000
	vk_structure_type_pipeline_viewport_swizzle_state_create_info_nv = 1000098000
	vk_structure_type_physical_device_discard_rectangle_properties_ext = 1000099000
	vk_structure_type_pipeline_discard_rectangle_state_create_info_ext = 1000099001
	vk_structure_type_physical_device_conservative_rasterization_properties_ext = 1000101000
	vk_structure_type_pipeline_rasterization_conservative_state_create_info_ext = 1000101001
	vk_structure_type_physical_device_depth_clip_enable_features_ext = 1000102000
	vk_structure_type_pipeline_rasterization_depth_clip_state_create_info_ext = 1000102001
	vk_structure_type_hdr_metadata_ext = 1000105000
	vk_structure_type_shared_present_surface_capabilities_khr = 1000111000
	vk_structure_type_import_fence_win32_handle_info_khr = 1000114000
	vk_structure_type_export_fence_win32_handle_info_khr = 1000114001
	vk_structure_type_fence_get_win32_handle_info_khr = 1000114002
	vk_structure_type_import_fence_fd_info_khr = 1000115000
	vk_structure_type_fence_get_fd_info_khr = 1000115001
	vk_structure_type_physical_device_performance_query_features_khr = 1000116000
	vk_structure_type_physical_device_performance_query_properties_khr = 1000116001
	vk_structure_type_query_pool_performance_create_info_khr = 1000116002
	vk_structure_type_performance_query_submit_info_khr = 1000116003
	vk_structure_type_acquire_profiling_lock_info_khr = 1000116004
	vk_structure_type_performance_counter_khr = 1000116005
	vk_structure_type_performance_counter_description_khr = 1000116006
	vk_structure_type_physical_device_surface_info_2_khr = 1000119000
	vk_structure_type_surface_capabilities_2_khr = 1000119001
	vk_structure_type_surface_format_2_khr = 1000119002
	vk_structure_type_display_properties_2_khr = 1000121000
	vk_structure_type_display_plane_properties_2_khr = 1000121001
	vk_structure_type_display_mode_properties_2_khr = 1000121002
	vk_structure_type_display_plane_info_2_khr = 1000121003
	vk_structure_type_display_plane_capabilities_2_khr = 1000121004
	vk_structure_type_ios_surface_create_info_mvk = 1000122000
	vk_structure_type_macos_surface_create_info_mvk = 1000123000
	vk_structure_type_debug_utils_object_name_info_ext = 1000128000
	vk_structure_type_debug_utils_object_tag_info_ext = 1000128001
	vk_structure_type_debug_utils_label_ext = 1000128002
	vk_structure_type_debug_utils_messenger_callback_data_ext = 1000128003
	vk_structure_type_debug_utils_messenger_create_info_ext = 1000128004
	vk_structure_type_android_hardware_buffer_usage_android = 1000129000
	vk_structure_type_android_hardware_buffer_properties_android = 1000129001
	vk_structure_type_android_hardware_buffer_format_properties_android = 1000129002
	vk_structure_type_import_android_hardware_buffer_info_android = 1000129003
	vk_structure_type_memory_get_android_hardware_buffer_info_android = 1000129004
	vk_structure_type_external_format_android = 1000129005
	vk_structure_type_physical_device_inline_uniform_block_features_ext = 1000138000
	vk_structure_type_physical_device_inline_uniform_block_properties_ext = 1000138001
	vk_structure_type_write_descriptor_set_inline_uniform_block_ext = 1000138002
	vk_structure_type_descriptor_pool_inline_uniform_block_create_info_ext = 1000138003
	vk_structure_type_sample_locations_info_ext = 1000143000
	vk_structure_type_render_pass_sample_locations_begin_info_ext = 1000143001
	vk_structure_type_pipeline_sample_locations_state_create_info_ext = 1000143002
	vk_structure_type_physical_device_sample_locations_properties_ext = 1000143003
	vk_structure_type_multisample_properties_ext = 1000143004
	vk_structure_type_physical_device_blend_operation_advanced_features_ext = 1000148000
	vk_structure_type_physical_device_blend_operation_advanced_properties_ext = 1000148001
	vk_structure_type_pipeline_color_blend_advanced_state_create_info_ext = 1000148002
	vk_structure_type_pipeline_coverage_to_color_state_create_info_nv = 1000149000
	vk_structure_type_write_descriptor_set_acceleration_structure_khr = 1000150007
	vk_structure_type_acceleration_structure_build_geometry_info_khr = 1000150000
	vk_structure_type_acceleration_structure_device_address_info_khr = 1000150002
	vk_structure_type_acceleration_structure_geometry_aabbs_data_khr = 1000150003
	vk_structure_type_acceleration_structure_geometry_instances_data_khr = 1000150004
	vk_structure_type_acceleration_structure_geometry_triangles_data_khr = 1000150005
	vk_structure_type_acceleration_structure_geometry_khr = 1000150006
	vk_structure_type_acceleration_structure_version_info_khr = 1000150009
	vk_structure_type_copy_acceleration_structure_info_khr = 1000150010
	vk_structure_type_copy_acceleration_structure_to_memory_info_khr = 1000150011
	vk_structure_type_copy_memory_to_acceleration_structure_info_khr = 1000150012
	vk_structure_type_physical_device_acceleration_structure_features_khr = 1000150013
	vk_structure_type_physical_device_acceleration_structure_properties_khr = 1000150014
	vk_structure_type_acceleration_structure_create_info_khr = 1000150017
	vk_structure_type_acceleration_structure_build_sizes_info_khr = 1000150020
	vk_structure_type_physical_device_ray_tracing_pipeline_features_khr = 1000347000
	vk_structure_type_physical_device_ray_tracing_pipeline_properties_khr = 1000347001
	vk_structure_type_ray_tracing_pipeline_create_info_khr = 1000150015
	vk_structure_type_ray_tracing_shader_group_create_info_khr = 1000150016
	vk_structure_type_ray_tracing_pipeline_interface_create_info_khr = 1000150018
	vk_structure_type_physical_device_ray_query_features_khr = 1000348013
	vk_structure_type_pipeline_coverage_modulation_state_create_info_nv = 1000152000
	vk_structure_type_physical_device_shader_sm_builtins_features_nv = 1000154000
	vk_structure_type_physical_device_shader_sm_builtins_properties_nv = 1000154001
	vk_structure_type_drm_format_modifier_properties_list_ext = 1000158000
	vk_structure_type_physical_device_image_drm_format_modifier_info_ext = 1000158002
	vk_structure_type_image_drm_format_modifier_list_create_info_ext = 1000158003
	vk_structure_type_image_drm_format_modifier_explicit_create_info_ext = 1000158004
	vk_structure_type_image_drm_format_modifier_properties_ext = 1000158005
	vk_structure_type_validation_cache_create_info_ext = 1000160000
	vk_structure_type_shader_module_validation_cache_create_info_ext = 1000160001
	vk_structure_type_physical_device_portability_subset_features_khr = 1000163000
	vk_structure_type_physical_device_portability_subset_properties_khr = 1000163001
	vk_structure_type_pipeline_viewport_shading_rate_image_state_create_info_nv = 1000164000
	vk_structure_type_physical_device_shading_rate_image_features_nv = 1000164001
	vk_structure_type_physical_device_shading_rate_image_properties_nv = 1000164002
	vk_structure_type_pipeline_viewport_coarse_sample_order_state_create_info_nv = 1000164005
	vk_structure_type_ray_tracing_pipeline_create_info_nv = 1000165000
	vk_structure_type_acceleration_structure_create_info_nv = 1000165001
	vk_structure_type_geometry_nv = 1000165003
	vk_structure_type_geometry_triangles_nv = 1000165004
	vk_structure_type_geometry_aabb_nv = 1000165005
	vk_structure_type_bind_acceleration_structure_memory_info_nv = 1000165006
	vk_structure_type_write_descriptor_set_acceleration_structure_nv = 1000165007
	vk_structure_type_acceleration_structure_memory_requirements_info_nv = 1000165008
	vk_structure_type_physical_device_ray_tracing_properties_nv = 1000165009
	vk_structure_type_ray_tracing_shader_group_create_info_nv = 1000165011
	vk_structure_type_acceleration_structure_info_nv = 1000165012
	vk_structure_type_physical_device_representative_fragment_test_features_nv = 1000166000
	vk_structure_type_pipeline_representative_fragment_test_state_create_info_nv = 1000166001
	vk_structure_type_physical_device_image_view_image_format_info_ext = 1000170000
	vk_structure_type_filter_cubic_image_view_image_format_properties_ext = 1000170001
	vk_structure_type_device_queue_global_priority_create_info_ext = 1000174000
	vk_structure_type_import_memory_host_pointer_info_ext = 1000178000
	vk_structure_type_memory_host_pointer_properties_ext = 1000178001
	vk_structure_type_physical_device_external_memory_host_properties_ext = 1000178002
	vk_structure_type_physical_device_shader_clock_features_khr = 1000181000
	vk_structure_type_pipeline_compiler_control_create_info_amd = 1000183000
	vk_structure_type_calibrated_timestamp_info_ext = 1000184000
	vk_structure_type_physical_device_shader_core_properties_amd = 1000185000
	vk_structure_type_video_decode_h265_capabilities_ext = 1000187000
	vk_structure_type_video_decode_h265_session_create_info_ext = 1000187001
	vk_structure_type_video_decode_h265_session_parameters_create_info_ext = 1000187002
	vk_structure_type_video_decode_h265_session_parameters_add_info_ext = 1000187003
	vk_structure_type_video_decode_h265_profile_ext = 1000187004
	vk_structure_type_video_decode_h265_picture_info_ext = 1000187005
	vk_structure_type_video_decode_h265_dpb_slot_info_ext = 1000187006
	vk_structure_type_device_memory_overallocation_create_info_amd = 1000189000
	vk_structure_type_physical_device_vertex_attribute_divisor_properties_ext = 1000190000
	vk_structure_type_pipeline_vertex_input_divisor_state_create_info_ext = 1000190001
	vk_structure_type_physical_device_vertex_attribute_divisor_features_ext = 1000190002
	vk_structure_type_present_frame_token_ggp = 1000191000
	vk_structure_type_pipeline_creation_feedback_create_info_ext = 1000192000
	vk_structure_type_physical_device_compute_shader_derivatives_features_nv = 1000201000
	vk_structure_type_physical_device_mesh_shader_features_nv = 1000202000
	vk_structure_type_physical_device_mesh_shader_properties_nv = 1000202001
	vk_structure_type_physical_device_fragment_shader_barycentric_features_nv = 1000203000
	vk_structure_type_physical_device_shader_image_footprint_features_nv = 1000204000
	vk_structure_type_pipeline_viewport_exclusive_scissor_state_create_info_nv = 1000205000
	vk_structure_type_physical_device_exclusive_scissor_features_nv = 1000205002
	vk_structure_type_checkpoint_data_nv = 1000206000
	vk_structure_type_queue_family_checkpoint_properties_nv = 1000206001
	vk_structure_type_physical_device_shader_integer_functions_2_features_intel = 1000209000
	vk_structure_type_query_pool_performance_query_create_info_intel = 1000210000
	vk_structure_type_initialize_performance_api_info_intel = 1000210001
	vk_structure_type_performance_marker_info_intel = 1000210002
	vk_structure_type_performance_stream_marker_info_intel = 1000210003
	vk_structure_type_performance_override_info_intel = 1000210004
	vk_structure_type_performance_configuration_acquire_info_intel = 1000210005
	vk_structure_type_physical_device_pci_bus_info_properties_ext = 1000212000
	vk_structure_type_display_native_hdr_surface_capabilities_amd = 1000213000
	vk_structure_type_swapchain_display_native_hdr_create_info_amd = 1000213001
	vk_structure_type_imagepipe_surface_create_info_fuchsia = 1000214000
	vk_structure_type_physical_device_shader_terminate_invocation_features_khr = 1000215000
	vk_structure_type_metal_surface_create_info_ext = 1000217000
	vk_structure_type_physical_device_fragment_density_map_features_ext = 1000218000
	vk_structure_type_physical_device_fragment_density_map_properties_ext = 1000218001
	vk_structure_type_render_pass_fragment_density_map_create_info_ext = 1000218002
	vk_structure_type_physical_device_subgroup_size_control_properties_ext = 1000225000
	vk_structure_type_pipeline_shader_stage_required_subgroup_size_create_info_ext = 1000225001
	vk_structure_type_physical_device_subgroup_size_control_features_ext = 1000225002
	vk_structure_type_fragment_shading_rate_attachment_info_khr = 1000226000
	vk_structure_type_pipeline_fragment_shading_rate_state_create_info_khr = 1000226001
	vk_structure_type_physical_device_fragment_shading_rate_properties_khr = 1000226002
	vk_structure_type_physical_device_fragment_shading_rate_features_khr = 1000226003
	vk_structure_type_physical_device_fragment_shading_rate_khr = 1000226004
	vk_structure_type_physical_device_shader_core_properties_2_amd = 1000227000
	vk_structure_type_physical_device_coherent_memory_features_amd = 1000229000
	vk_structure_type_physical_device_shader_image_atomic_int64_features_ext = 1000234000
	vk_structure_type_physical_device_memory_budget_properties_ext = 1000237000
	vk_structure_type_physical_device_memory_priority_features_ext = 1000238000
	vk_structure_type_memory_priority_allocate_info_ext = 1000238001
	vk_structure_type_surface_protected_capabilities_khr = 1000239000
	vk_structure_type_physical_device_dedicated_allocation_image_aliasing_features_nv = 1000240000
	vk_structure_type_physical_device_buffer_device_address_features_ext = 1000244000
	vk_structure_type_buffer_device_address_create_info_ext = 1000244002
	vk_structure_type_physical_device_tool_properties_ext = 1000245000
	vk_structure_type_validation_features_ext = 1000247000
	vk_structure_type_physical_device_present_wait_features_khr = 1000248000
	vk_structure_type_physical_device_cooperative_matrix_features_nv = 1000249000
	vk_structure_type_cooperative_matrix_properties_nv = 1000249001
	vk_structure_type_physical_device_cooperative_matrix_properties_nv = 1000249002
	vk_structure_type_physical_device_coverage_reduction_mode_features_nv = 1000250000
	vk_structure_type_pipeline_coverage_reduction_state_create_info_nv = 1000250001
	vk_structure_type_framebuffer_mixed_samples_combination_nv = 1000250002
	vk_structure_type_physical_device_fragment_shader_interlock_features_ext = 1000251000
	vk_structure_type_physical_device_ycbcr_image_arrays_features_ext = 1000252000
	vk_structure_type_physical_device_provoking_vertex_features_ext = 1000254000
	vk_structure_type_pipeline_rasterization_provoking_vertex_state_create_info_ext = 1000254001
	vk_structure_type_physical_device_provoking_vertex_properties_ext = 1000254002
	vk_structure_type_surface_full_screen_exclusive_info_ext = 1000255000
	vk_structure_type_surface_capabilities_full_screen_exclusive_ext = 1000255002
	vk_structure_type_surface_full_screen_exclusive_win32_info_ext = 1000255001
	vk_structure_type_headless_surface_create_info_ext = 1000256000
	vk_structure_type_physical_device_line_rasterization_features_ext = 1000259000
	vk_structure_type_pipeline_rasterization_line_state_create_info_ext = 1000259001
	vk_structure_type_physical_device_line_rasterization_properties_ext = 1000259002
	vk_structure_type_physical_device_shader_atomic_float_features_ext = 1000260000
	vk_structure_type_physical_device_index_type_uint8_features_ext = 1000265000
	vk_structure_type_physical_device_extended_dynamic_state_features_ext = 1000267000
	vk_structure_type_physical_device_pipeline_executable_properties_features_khr = 1000269000
	vk_structure_type_pipeline_info_khr = 1000269001
	vk_structure_type_pipeline_executable_properties_khr = 1000269002
	vk_structure_type_pipeline_executable_info_khr = 1000269003
	vk_structure_type_pipeline_executable_statistic_khr = 1000269004
	vk_structure_type_pipeline_executable_internal_representation_khr = 1000269005
	vk_structure_type_physical_device_shader_atomic_float_2_features_ext = 1000273000
	vk_structure_type_physical_device_shader_demote_to_helper_invocation_features_ext = 1000276000
	vk_structure_type_physical_device_device_generated_commands_properties_nv = 1000277000
	vk_structure_type_graphics_shader_group_create_info_nv = 1000277001
	vk_structure_type_graphics_pipeline_shader_groups_create_info_nv = 1000277002
	vk_structure_type_indirect_commands_layout_token_nv = 1000277003
	vk_structure_type_indirect_commands_layout_create_info_nv = 1000277004
	vk_structure_type_generated_commands_info_nv = 1000277005
	vk_structure_type_generated_commands_memory_requirements_info_nv = 1000277006
	vk_structure_type_physical_device_device_generated_commands_features_nv = 1000277007
	vk_structure_type_physical_device_inherited_viewport_scissor_features_nv = 1000278000
	vk_structure_type_command_buffer_inheritance_viewport_scissor_info_nv = 1000278001
	vk_structure_type_physical_device_texel_buffer_alignment_features_ext = 1000281000
	vk_structure_type_physical_device_texel_buffer_alignment_properties_ext = 1000281001
	vk_structure_type_command_buffer_inheritance_render_pass_transform_info_qcom = 1000282000
	vk_structure_type_render_pass_transform_begin_info_qcom = 1000282001
	vk_structure_type_physical_device_device_memory_report_features_ext = 1000284000
	vk_structure_type_device_device_memory_report_create_info_ext = 1000284001
	vk_structure_type_device_memory_report_callback_data_ext = 1000284002
	vk_structure_type_physical_device_robustness_2_features_ext = 1000286000
	vk_structure_type_physical_device_robustness_2_properties_ext = 1000286001
	vk_structure_type_sampler_custom_border_color_create_info_ext = 1000287000
	vk_structure_type_physical_device_custom_border_color_properties_ext = 1000287001
	vk_structure_type_physical_device_custom_border_color_features_ext = 1000287002
	vk_structure_type_pipeline_library_create_info_khr = 1000290000
	vk_structure_type_present_id_khr = 1000294000
	vk_structure_type_physical_device_present_id_features_khr = 1000294001
	vk_structure_type_physical_device_private_data_features_ext = 1000295000
	vk_structure_type_device_private_data_create_info_ext = 1000295001
	vk_structure_type_private_data_slot_create_info_ext = 1000295002
	vk_structure_type_physical_device_pipeline_creation_cache_control_features_ext = 1000297000
	vk_structure_type_video_encode_info_khr = 1000299000
	vk_structure_type_video_encode_rate_control_info_khr = 1000299001
	vk_structure_type_physical_device_diagnostics_config_features_nv = 1000300000
	vk_structure_type_device_diagnostics_config_create_info_nv = 1000300001
	vk_structure_type_memory_barrier_2_khr = 1000314000
	vk_structure_type_buffer_memory_barrier_2_khr = 1000314001
	vk_structure_type_image_memory_barrier_2_khr = 1000314002
	vk_structure_type_dependency_info_khr = 1000314003
	vk_structure_type_submit_info_2_khr = 1000314004
	vk_structure_type_semaphore_submit_info_khr = 1000314005
	vk_structure_type_command_buffer_submit_info_khr = 1000314006
	vk_structure_type_physical_device_synchronization_2_features_khr = 1000314007
	vk_structure_type_queue_family_checkpoint_properties_2_nv = 1000314008
	vk_structure_type_checkpoint_data_2_nv = 1000314009
	vk_structure_type_physical_device_shader_subgroup_uniform_control_flow_features_khr = 1000323000
	vk_structure_type_physical_device_zero_initialize_workgroup_memory_features_khr = 1000325000
	vk_structure_type_physical_device_fragment_shading_rate_enums_properties_nv = 1000326000
	vk_structure_type_physical_device_fragment_shading_rate_enums_features_nv = 1000326001
	vk_structure_type_pipeline_fragment_shading_rate_enum_state_create_info_nv = 1000326002
	vk_structure_type_acceleration_structure_geometry_motion_triangles_data_nv = 1000327000
	vk_structure_type_physical_device_ray_tracing_motion_blur_features_nv = 1000327001
	vk_structure_type_acceleration_structure_motion_info_nv = 1000327002
	vk_structure_type_physical_device_ycbcr_2_plane_444_formats_features_ext = 1000330000
	vk_structure_type_physical_device_fragment_density_map_2_features_ext = 1000332000
	vk_structure_type_physical_device_fragment_density_map_2_properties_ext = 1000332001
	vk_structure_type_copy_command_transform_info_qcom = 1000333000
	vk_structure_type_physical_device_image_robustness_features_ext = 1000335000
	vk_structure_type_physical_device_workgroup_memory_explicit_layout_features_khr = 1000336000
	vk_structure_type_copy_buffer_info_2_khr = 1000337000
	vk_structure_type_copy_image_info_2_khr = 1000337001
	vk_structure_type_copy_buffer_to_image_info_2_khr = 1000337002
	vk_structure_type_copy_image_to_buffer_info_2_khr = 1000337003
	vk_structure_type_blit_image_info_2_khr = 1000337004
	vk_structure_type_resolve_image_info_2_khr = 1000337005
	vk_structure_type_buffer_copy_2_khr = 1000337006
	vk_structure_type_image_copy_2_khr = 1000337007
	vk_structure_type_image_blit_2_khr = 1000337008
	vk_structure_type_buffer_image_copy_2_khr = 1000337009
	vk_structure_type_image_resolve_2_khr = 1000337010
	vk_structure_type_physical_device_4444_formats_features_ext = 1000340000
	vk_structure_type_directfb_surface_create_info_ext = 1000346000
	vk_structure_type_physical_device_mutable_descriptor_type_features_valve = 1000351000
	vk_structure_type_mutable_descriptor_type_create_info_valve = 1000351002
	vk_structure_type_physical_device_vertex_input_dynamic_state_features_ext = 1000352000
	vk_structure_type_vertex_input_binding_description_2_ext = 1000352001
	vk_structure_type_vertex_input_attribute_description_2_ext = 1000352002
	vk_structure_type_physical_device_drm_properties_ext = 1000353000
	vk_structure_type_import_memory_zircon_handle_info_fuchsia = 1000364000
	vk_structure_type_memory_zircon_handle_properties_fuchsia = 1000364001
	vk_structure_type_memory_get_zircon_handle_info_fuchsia = 1000364002
	vk_structure_type_import_semaphore_zircon_handle_info_fuchsia = 1000365000
	vk_structure_type_semaphore_get_zircon_handle_info_fuchsia = 1000365001
	vk_structure_type_subpass_shading_pipeline_create_info_huawei = 1000369000
	vk_structure_type_physical_device_subpass_shading_features_huawei = 1000369001
	vk_structure_type_physical_device_subpass_shading_properties_huawei = 1000369002
	vk_structure_type_physical_device_invocation_mask_features_huawei = 1000370000
	vk_structure_type_memory_get_remote_address_info_nv = 1000371000
	vk_structure_type_physical_device_external_memory_rdma_features_nv = 1000371001
	vk_structure_type_physical_device_extended_dynamic_state_2_features_ext = 1000377000
	vk_structure_type_screen_surface_create_info_qnx = 1000378000
	vk_structure_type_physical_device_color_write_enable_features_ext = 1000381000
	vk_structure_type_pipeline_color_write_create_info_ext = 1000381001
	vk_structure_type_physical_device_global_priority_query_features_ext = 1000388000
	vk_structure_type_queue_family_global_priority_properties_ext = 1000388001
	vk_structure_type_physical_device_multi_draw_features_ext = 1000392000
	vk_structure_type_physical_device_multi_draw_properties_ext = 1000392001
	/*
	vk_structure_type_physical_device_variable_pointer_features = vk_structure_type_physical_device_variable_pointers_features
	vk_structure_type_physical_device_shader_draw_parameter_features = vk_structure_type_physical_device_shader_draw_parameters_features
	vk_structure_type_debug_report_create_info_ext = vk_structure_type_debug_report_callback_create_info_ext
	vk_structure_type_render_pass_multiview_create_info_khr = vk_structure_type_render_pass_multiview_create_info
	vk_structure_type_physical_device_multiview_features_khr = vk_structure_type_physical_device_multiview_features
	vk_structure_type_physical_device_multiview_properties_khr = vk_structure_type_physical_device_multiview_properties
	vk_structure_type_physical_device_features_2_khr = vk_structure_type_physical_device_features_2
	vk_structure_type_physical_device_properties_2_khr = vk_structure_type_physical_device_properties_2
	vk_structure_type_format_properties_2_khr = vk_structure_type_format_properties_2
	vk_structure_type_image_format_properties_2_khr = vk_structure_type_image_format_properties_2
	vk_structure_type_physical_device_image_format_info_2_khr = vk_structure_type_physical_device_image_format_info_2
	vk_structure_type_queue_family_properties_2_khr = vk_structure_type_queue_family_properties_2
	vk_structure_type_physical_device_memory_properties_2_khr = vk_structure_type_physical_device_memory_properties_2
	vk_structure_type_sparse_image_format_properties_2_khr = vk_structure_type_sparse_image_format_properties_2
	vk_structure_type_physical_device_sparse_image_format_info_2_khr = vk_structure_type_physical_device_sparse_image_format_info_2
	vk_structure_type_memory_allocate_flags_info_khr = vk_structure_type_memory_allocate_flags_info
	vk_structure_type_device_group_render_pass_begin_info_khr = vk_structure_type_device_group_render_pass_begin_info
	vk_structure_type_device_group_command_buffer_begin_info_khr = vk_structure_type_device_group_command_buffer_begin_info
	vk_structure_type_device_group_submit_info_khr = vk_structure_type_device_group_submit_info
	vk_structure_type_device_group_bind_sparse_info_khr = vk_structure_type_device_group_bind_sparse_info
	vk_structure_type_bind_buffer_memory_device_group_info_khr = vk_structure_type_bind_buffer_memory_device_group_info
	vk_structure_type_bind_image_memory_device_group_info_khr = vk_structure_type_bind_image_memory_device_group_info
	vk_structure_type_physical_device_group_properties_khr = vk_structure_type_physical_device_group_properties
	vk_structure_type_device_group_device_create_info_khr = vk_structure_type_device_group_device_create_info
	vk_structure_type_physical_device_external_image_format_info_khr = vk_structure_type_physical_device_external_image_format_info
	vk_structure_type_external_image_format_properties_khr = vk_structure_type_external_image_format_properties
	vk_structure_type_physical_device_external_buffer_info_khr = vk_structure_type_physical_device_external_buffer_info
	vk_structure_type_external_buffer_properties_khr = vk_structure_type_external_buffer_properties
	vk_structure_type_physical_device_id_properties_khr = vk_structure_type_physical_device_id_properties
	vk_structure_type_external_memory_buffer_create_info_khr = vk_structure_type_external_memory_buffer_create_info
	vk_structure_type_external_memory_image_create_info_khr = vk_structure_type_external_memory_image_create_info
	vk_structure_type_export_memory_allocate_info_khr = vk_structure_type_export_memory_allocate_info
	vk_structure_type_physical_device_external_semaphore_info_khr = vk_structure_type_physical_device_external_semaphore_info
	vk_structure_type_external_semaphore_properties_khr = vk_structure_type_external_semaphore_properties
	vk_structure_type_export_semaphore_create_info_khr = vk_structure_type_export_semaphore_create_info
	vk_structure_type_physical_device_shader_float16_int8_features_khr = vk_structure_type_physical_device_shader_float16_int8_features
	vk_structure_type_physical_device_float16_int8_features_khr = vk_structure_type_physical_device_shader_float16_int8_features
	vk_structure_type_physical_device_16bit_storage_features_khr = vk_structure_type_physical_device_16bit_storage_features
	vk_structure_type_descriptor_update_template_create_info_khr = vk_structure_type_descriptor_update_template_create_info
	vk_structure_type_surface_capabilities2_ext = vk_structure_type_surface_capabilities_2_ext
	vk_structure_type_physical_device_imageless_framebuffer_features_khr = vk_structure_type_physical_device_imageless_framebuffer_features
	vk_structure_type_framebuffer_attachments_create_info_khr = vk_structure_type_framebuffer_attachments_create_info
	vk_structure_type_framebuffer_attachment_image_info_khr = vk_structure_type_framebuffer_attachment_image_info
	vk_structure_type_render_pass_attachment_begin_info_khr = vk_structure_type_render_pass_attachment_begin_info
	vk_structure_type_attachment_description_2_khr = vk_structure_type_attachment_description_2
	vk_structure_type_attachment_reference_2_khr = vk_structure_type_attachment_reference_2
	vk_structure_type_subpass_description_2_khr = vk_structure_type_subpass_description_2
	vk_structure_type_subpass_dependency_2_khr = vk_structure_type_subpass_dependency_2
	vk_structure_type_render_pass_create_info_2_khr = vk_structure_type_render_pass_create_info_2
	vk_structure_type_subpass_begin_info_khr = vk_structure_type_subpass_begin_info
	vk_structure_type_subpass_end_info_khr = vk_structure_type_subpass_end_info
	vk_structure_type_physical_device_external_fence_info_khr = vk_structure_type_physical_device_external_fence_info
	vk_structure_type_external_fence_properties_khr = vk_structure_type_external_fence_properties
	vk_structure_type_export_fence_create_info_khr = vk_structure_type_export_fence_create_info
	vk_structure_type_physical_device_point_clipping_properties_khr = vk_structure_type_physical_device_point_clipping_properties
	vk_structure_type_render_pass_input_attachment_aspect_create_info_khr = vk_structure_type_render_pass_input_attachment_aspect_create_info
	vk_structure_type_image_view_usage_create_info_khr = vk_structure_type_image_view_usage_create_info
	vk_structure_type_pipeline_tessellation_domain_origin_state_create_info_khr = vk_structure_type_pipeline_tessellation_domain_origin_state_create_info
	vk_structure_type_physical_device_variable_pointers_features_khr = vk_structure_type_physical_device_variable_pointers_features
	vk_structure_type_physical_device_variable_pointer_features_khr = vk_structure_type_physical_device_variable_pointers_features_khr
	vk_structure_type_memory_dedicated_requirements_khr = vk_structure_type_memory_dedicated_requirements
	vk_structure_type_memory_dedicated_allocate_info_khr = vk_structure_type_memory_dedicated_allocate_info
	vk_structure_type_physical_device_sampler_filter_minmax_properties_ext = vk_structure_type_physical_device_sampler_filter_minmax_properties
	vk_structure_type_sampler_reduction_mode_create_info_ext = vk_structure_type_sampler_reduction_mode_create_info
	vk_structure_type_buffer_memory_requirements_info_2_khr = vk_structure_type_buffer_memory_requirements_info_2
	vk_structure_type_image_memory_requirements_info_2_khr = vk_structure_type_image_memory_requirements_info_2
	vk_structure_type_image_sparse_memory_requirements_info_2_khr = vk_structure_type_image_sparse_memory_requirements_info_2
	vk_structure_type_memory_requirements_2_khr = vk_structure_type_memory_requirements_2
	vk_structure_type_sparse_image_memory_requirements_2_khr = vk_structure_type_sparse_image_memory_requirements_2
	vk_structure_type_image_format_list_create_info_khr = vk_structure_type_image_format_list_create_info
	vk_structure_type_sampler_ycbcr_conversion_create_info_khr = vk_structure_type_sampler_ycbcr_conversion_create_info
	vk_structure_type_sampler_ycbcr_conversion_info_khr = vk_structure_type_sampler_ycbcr_conversion_info
	vk_structure_type_bind_image_plane_memory_info_khr = vk_structure_type_bind_image_plane_memory_info
	vk_structure_type_image_plane_memory_requirements_info_khr = vk_structure_type_image_plane_memory_requirements_info
	vk_structure_type_physical_device_sampler_ycbcr_conversion_features_khr = vk_structure_type_physical_device_sampler_ycbcr_conversion_features
	vk_structure_type_sampler_ycbcr_conversion_image_format_properties_khr = vk_structure_type_sampler_ycbcr_conversion_image_format_properties
	vk_structure_type_bind_buffer_memory_info_khr = vk_structure_type_bind_buffer_memory_info
	vk_structure_type_bind_image_memory_info_khr = vk_structure_type_bind_image_memory_info
	vk_structure_type_descriptor_set_layout_binding_flags_create_info_ext = vk_structure_type_descriptor_set_layout_binding_flags_create_info
	vk_structure_type_physical_device_descriptor_indexing_features_ext = vk_structure_type_physical_device_descriptor_indexing_features
	vk_structure_type_physical_device_descriptor_indexing_properties_ext = vk_structure_type_physical_device_descriptor_indexing_properties
	vk_structure_type_descriptor_set_variable_descriptor_count_allocate_info_ext = vk_structure_type_descriptor_set_variable_descriptor_count_allocate_info
	vk_structure_type_descriptor_set_variable_descriptor_count_layout_support_ext = vk_structure_type_descriptor_set_variable_descriptor_count_layout_support
	vk_structure_type_physical_device_maintenance_3_properties_khr = vk_structure_type_physical_device_maintenance_3_properties
	vk_structure_type_descriptor_set_layout_support_khr = vk_structure_type_descriptor_set_layout_support
	vk_structure_type_physical_device_shader_subgroup_extended_types_features_khr = vk_structure_type_physical_device_shader_subgroup_extended_types_features
	vk_structure_type_physical_device_8bit_storage_features_khr = vk_structure_type_physical_device_8bit_storage_features
	vk_structure_type_physical_device_shader_atomic_int64_features_khr = vk_structure_type_physical_device_shader_atomic_int64_features
	vk_structure_type_physical_device_driver_properties_khr = vk_structure_type_physical_device_driver_properties
	vk_structure_type_physical_device_float_controls_properties_khr = vk_structure_type_physical_device_float_controls_properties
	vk_structure_type_physical_device_depth_stencil_resolve_properties_khr = vk_structure_type_physical_device_depth_stencil_resolve_properties
	vk_structure_type_subpass_description_depth_stencil_resolve_khr = vk_structure_type_subpass_description_depth_stencil_resolve
	vk_structure_type_physical_device_timeline_semaphore_features_khr = vk_structure_type_physical_device_timeline_semaphore_features
	vk_structure_type_physical_device_timeline_semaphore_properties_khr = vk_structure_type_physical_device_timeline_semaphore_properties
	vk_structure_type_semaphore_type_create_info_khr = vk_structure_type_semaphore_type_create_info
	vk_structure_type_timeline_semaphore_submit_info_khr = vk_structure_type_timeline_semaphore_submit_info
	vk_structure_type_semaphore_wait_info_khr = vk_structure_type_semaphore_wait_info
	vk_structure_type_semaphore_signal_info_khr = vk_structure_type_semaphore_signal_info
	vk_structure_type_query_pool_create_info_intel = vk_structure_type_query_pool_performance_query_create_info_intel
	vk_structure_type_physical_device_vulkan_memory_model_features_khr = vk_structure_type_physical_device_vulkan_memory_model_features
	vk_structure_type_physical_device_scalar_block_layout_features_ext = vk_structure_type_physical_device_scalar_block_layout_features
	vk_structure_type_physical_device_separate_depth_stencil_layouts_features_khr = vk_structure_type_physical_device_separate_depth_stencil_layouts_features
	vk_structure_type_attachment_reference_stencil_layout_khr = vk_structure_type_attachment_reference_stencil_layout
	vk_structure_type_attachment_description_stencil_layout_khr = vk_structure_type_attachment_description_stencil_layout
	vk_structure_type_physical_device_buffer_address_features_ext = vk_structure_type_physical_device_buffer_device_address_features_ext
	vk_structure_type_buffer_device_address_info_ext = vk_structure_type_buffer_device_address_info
	vk_structure_type_image_stencil_usage_create_info_ext = vk_structure_type_image_stencil_usage_create_info
	vk_structure_type_physical_device_uniform_buffer_standard_layout_features_khr = vk_structure_type_physical_device_uniform_buffer_standard_layout_features
	vk_structure_type_physical_device_buffer_device_address_features_khr = vk_structure_type_physical_device_buffer_device_address_features
	vk_structure_type_buffer_device_address_info_khr = vk_structure_type_buffer_device_address_info
	vk_structure_type_buffer_opaque_capture_address_create_info_khr = vk_structure_type_buffer_opaque_capture_address_create_info
	vk_structure_type_memory_opaque_capture_address_allocate_info_khr = vk_structure_type_memory_opaque_capture_address_allocate_info
	vk_structure_type_device_memory_opaque_capture_address_info_khr = vk_structure_type_device_memory_opaque_capture_address_info
	vk_structure_type_physical_device_host_query_reset_features_ext = vk_structure_type_physical_device_host_query_reset_features
	*/
	vk_structure_type_max_enum = 0x7fffffff
}
