module vulkan

#pkgconfig vulkan
#include <vulkan/vulkan.h>
