module vulkan

[heap; typedef]
struct C.VkSampleMask {}

[typedef]
struct C.VkPipelineLayout {}

[typedef]
struct C.VkDescriptorSetLayout {}

[typedef]
struct C.VkImageView {}

[typedef]
struct C.VkShaderModule {}

[typedef]
struct C.VkSwapchainKHR {}

[typedef]
struct C.VkBool32 {}

[typedef]
struct C.VkImage {}

[typedef]
struct C.VkDevice {}

[typedef]
struct C.VkQueue {}

[typedef]
struct C.VkSurfaceKHR {}

[typedef]
struct C.VkInstance {}

[typedef]
struct C.VkPhysicalDevice {}

[typedef]
struct C.VkRenderPass {}

[typedef]
struct C.VkPipeline {}

[typedef]
struct C.VkFramebuffer {}

[typedef]
struct C.VkCommandPool {}

[typedef]
struct C.VkCommandBuffer {}

[typedef]
struct C.VkSemaphore {}

[typedef]
struct C.VkFence {}

[typedef]
struct C.VkBuffer {}

[typedef]
struct C.VkDeviceMemory {}

[typedef]
struct C.VkDescriptorSetLayout {}

[typedef]
struct C.VkDescriptorPool {}

[typedef]
struct C.VkDescriptorSet {}

// TODO complete
[heap; typedef]
struct C.VkPipelineTessellationStateCreateInfo {}

[heap; typedef]
struct C.VkPipelineDepthStencilStateCreateInfo {}

[heap; typedef]
struct C.VkCommandBufferInheritanceInfo {}

[typedef]
struct C.VkPipelineCache {}

[typedef]
struct C.VkSampler {}
