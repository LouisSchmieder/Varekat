module mathf
